`include "parametersSiFH.vh"

module 4stateSiFH (
    ports
);
    
endmodule