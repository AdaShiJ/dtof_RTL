`include "parametersSiFH.vh"

module  algebraicBlock(
    input [`Nb:1] peakCH,
    //input peakReady,
    output reg [`Nb:1] THminus,
    output reg [`Nb:1] THpositive,
    output reg [`Nb:1] delta
);

reg [`Np:1] TTHminus;
reg [`Np:1] TTHpositive;
reg [`Np:1] SB;
reg [`Np:1] CH;
reg [`Np:1] upperBound;
reg [`Nb:1] upperBoundCH;

always @(*) begin
    upperBound <= ~0;
    upperBoundCH <= ~0;
    SB = 1 << (`Nb - 1); //32
    CH = peakCH << (`Np - `Nb);
    TTHminus = CH - SB;//bound
    TTHpositive = CH + SB;//bound
    if (CH >=  (upperBound - SB)) begin
        TTHpositive = upperBound - upperBoundCH;//wtf
        TTHminus = TTHpositive - 2* SB;
    end
    else begin
        if (CH <=  SB) begin
            TTHminus = 0;
            TTHpositive = TTHminus + 2* SB;
        end
        else begin
            TTHpositive = CH + SB;//wtf
            TTHminus = CH - SB;
        end
    end

    THminus <= TTHminus[`Np:`Np-`Nb+1];
    THpositive <= TTHpositive[`Np:`Np-`Nb+1];
    delta <= THminus + THpositive - (THpositive >> `Nb) << `Nb ;
end
    
endmodule