`include "parametersSiFH.vh"

module SiFHtop (
    ports
);
    
endmodule