`include "parametersSiFH.vh"

module  (
    ports 
);
    
endmodule