`define Nb 6
`define Np 10
`define peakMax 21
//`define peakMaxb = 15
//`define peakMaxp = 11