`define Nb 6
`define Np 10
`define NumberOfBins 64
`define peakMax 21
`define ACQ_NUM 4
`define DATA_NUM 2
`define SRAM_NUM 2
`define PIXEL_NUM 6
`define PIXEL_PER_RAM `PIXEL_NUM + `SRAM_NUM
`define RAM_SIZE `peakMax + `NUM_PER_RAM
`define ACQ_NUM_PER_RAM `ACQ_NUM + `PIXEL_PER_RAM

