`include "parametersSiFH.vh"

module topFSM (
    ports
);
    
endmodule