`define Nb 6
`define Np 10
`define NumberOfBins 64//2^(Nb)
`define peakMax 21
`define num_acq 4//33333
//`define peakMaxb = 15
//`define peakMaxp = 11