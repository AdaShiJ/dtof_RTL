`include "parametersSiFH.vh"

module peakDetecter (
    ports
);
    
endmodule


